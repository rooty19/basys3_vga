invader_tableTEMP[0]     <= 52'h0_000_000_20_0_ff0;
invader_tableTEMP[1]     <= 52'h0_000_020_20_0_ff0;
invader_tableTEMP[2]     <= 52'h0_000_040_20_0_ff0;
invader_tableTEMP[3]     <= 52'h0_000_060_20_0_ff0;
invader_tableTEMP[4]     <= 52'h0_000_0a0_20_0_ff0;
invader_tableTEMP[5]     <= 52'h0_000_0c0_20_0_ff0;
invader_tableTEMP[6]     <= 52'h0_000_0e0_20_0_ff0;
invader_tableTEMP[7]     <= 52'h0_000_100_20_0_ff0;
invader_tableTEMP[8]     <= 52'h0_030_000_20_0_0ff;
invader_tableTEMP[9]     <= 52'h0_030_020_20_0_0ff;
invader_tableTEMP[10]    <= 52'h0_030_040_20_0_0ff;
invader_tableTEMP[11]    <= 52'h0_030_060_20_0_0ff;
invader_tableTEMP[12]    <= 52'h0_030_0a0_20_0_0ff;
invader_tableTEMP[13]    <= 52'h0_030_0c0_20_0_0ff;
invader_tableTEMP[14]    <= 52'h0_030_0e0_20_0_0ff;
invader_tableTEMP[15]    <= 52'h0_030_100_20_0_0ff;
invader_tableTEMP[16]    <= 52'h0_060_000_20_0_f0f;
invader_tableTEMP[17]    <= 52'h0_060_020_20_0_f0f;
invader_tableTEMP[18]    <= 52'h0_060_040_20_0_f0f;
invader_tableTEMP[19]    <= 52'h0_060_060_20_0_f0f;
invader_tableTEMP[20]    <= 52'h0_060_0a0_20_0_f0f;
invader_tableTEMP[21]    <= 52'h0_060_0c0_20_0_f0f;
invader_tableTEMP[22]    <= 52'h0_060_0e0_20_0_f0f;
invader_tableTEMP[23]    <= 52'h0_060_100_20_0_f0f;
invader_tableTEMP[24]    <= 52'h0_090_000_20_0_fff;
invader_tableTEMP[25]    <= 52'h0_090_020_20_0_fff;
invader_tableTEMP[26]    <= 52'h0_090_040_20_0_fff;
invader_tableTEMP[27]    <= 52'h0_090_060_20_0_fff;
invader_tableTEMP[28]    <= 52'h0_090_0a0_20_0_fff;
invader_tableTEMP[29]    <= 52'h0_090_0c0_20_0_fff;
invader_tableTEMP[30]    <= 52'h0_090_0e0_20_0_fff;
invader_tableTEMP[31]    <= 52'h0_090_100_20_0_fff;
invader_tableTEMP[32]    <= 52'h0_020_1a0_20_0_fff;
invader_tableTEMP[33]    <= 52'h0_020_1c0_20_0_fff;
invader_tableTEMP[34]    <= 52'h0_020_1e0_20_0_fff;
invader_tableTEMP[35]    <= 52'h0_020_200_20_0_fff;
invader_tableTEMP[36]    <= 52'h0_020_220_20_0_fff;
invader_tableTEMP[37]    <= 52'h0_020_240_20_0_fff;
invader_tableTEMP[38]    <= 52'h0_020_260_20_0_fff;
invader_tableTEMP[39]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[40]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[41]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[42]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[43]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[44]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[45]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[46]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[47]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[48]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[50]    <= 52'h0_1c0_000_20_1_fff;
invader_tableTEMP[51]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[52]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[53]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[54]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[55]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[56]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[57]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[58]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[59]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[60]    <= 52'h0_000_000_20_0_000;
invader_tableTEMP[61]    <= 52'h0_1a0_000_20_1_000;
invader_tableTEMP[62]    <= 52'h0_1c0_000_20_1_ff0;