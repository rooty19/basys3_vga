            laser_table[0]  <= 40'h0_000_001_fff;
            laser_table[1]  <= 40'h0_000_010_ff0;
            laser_table[2]  <= 40'h0_000_000_000;
            laser_table[3]  <= 40'h0_000_000_000;
            laser_table[4]  <= 40'h0_000_000_000;
            laser_table[5]  <= 40'h0_000_000_000;
            laser_table[6]  <= 40'h0_000_000_000;
            laser_table[7]  <= 40'h0_000_000_000;
            laser_table[8]  <= 40'h0_000_000_000;
            laser_table[9]  <= 40'h0_000_020_ff0;
            laser_table[10] <= 40'h0_000_000_000;
            laser_table[11]  <= 40'h0_000_000_000;
            laser_table[12]  <= 40'h0_000_000_000;
            laser_table[13]  <= 40'h0_000_030_ff0;
            laser_table[14]  <= 40'h0_000_000_000;
            laser_table[15]  <= 40'h0_000_000_000;
            laser_table[16]  <= 40'h0_000_000_000;
            laser_table[17]  <= 40'h0_000_000_000;
            laser_table[18]  <= 40'h0_000_000_000;
            laser_table[19]  <= 40'h0_000_040_ff0;
            laser_table[20]  <= 40'h0_000_000_000;
            laser_table[21]  <= 40'h0_000_000_000;
            laser_table[22]  <= 40'h0_000_000_000;
            laser_table[23]  <= 40'h0_000_000_000;
            laser_table[24]  <= 40'h0_000_000_000;
            laser_table[25]  <= 40'h0_000_050_ff0;
            laser_table[26]  <= 40'h0_000_000_000;
            laser_table[27]  <= 40'h0_000_000_000;
            laser_table[28]  <= 40'h0_000_000_000;
            laser_table[29]  <= 40'h0_000_000_000;
            laser_table[30]  <= 40'h0_000_060_ff0;
            laser_table[31]  <= 40'h0_000_000_000;
            laser_table[32]  <= 40'h0_000_000_000;
            laser_table[33]  <= 40'h0_000_000_000;
            laser_table[34]  <= 40'h0_000_000_000;
            laser_table[35]  <= 40'h0_000_000_000;
            laser_table[36]  <= 40'h0_000_070_ff0;
            laser_table[37]  <= 40'h0_000_000_000;
            laser_table[38]  <= 40'h0_000_000_000;
            laser_table[39]  <= 40'h0_000_080_ff0;