invader_table[0]     <= 52'h8_000_000_20_0_ff0;
invader_table[1]     <= 52'h8_000_020_20_0_ff0;
invader_table[2]     <= 52'h8_000_040_20_0_ff0;
invader_table[3]     <= 52'h8_000_060_20_0_ff0;
invader_table[4]     <= 52'h8_000_0a0_20_0_ff0;
invader_table[5]     <= 52'h8_000_0c0_20_0_ff0;
invader_table[6]     <= 52'h8_000_0e0_20_0_ff0;
invader_table[7]     <= 52'h8_000_100_20_0_ff0;
invader_table[8]     <= 52'h8_030_000_20_0_0ff;
invader_table[9]     <= 52'h8_030_020_20_0_0ff;
invader_table[10]    <= 52'h8_030_040_20_0_0ff;
invader_table[11]    <= 52'h8_030_060_20_0_0ff;
invader_table[12]    <= 52'h8_030_0a0_20_0_0ff;
invader_table[13]    <= 52'h8_030_0c0_20_0_0ff;
invader_table[14]    <= 52'h8_030_0e0_20_0_0ff;
invader_table[15]    <= 52'h8_030_100_20_0_0ff;
invader_table[16]    <= 52'h8_060_000_20_0_f0f;
invader_table[17]    <= 52'h8_060_020_20_0_f0f;
invader_table[18]    <= 52'h8_060_040_20_0_f0f;
invader_table[19]    <= 52'h8_060_060_20_0_f0f;
invader_table[20]    <= 52'h8_060_0a0_20_0_f0f;
invader_table[21]    <= 52'h8_060_0c0_20_0_f0f;
invader_table[22]    <= 52'h8_060_0e0_20_0_f0f;
invader_table[23]    <= 52'h8_060_100_20_0_f0f;
invader_table[24]    <= 52'h8_090_000_20_0_fff;
invader_table[25]    <= 52'h8_090_020_20_0_fff;
invader_table[26]    <= 52'h8_090_040_20_0_fff;
invader_table[27]    <= 52'h8_090_060_20_0_fff;
invader_table[28]    <= 52'h8_090_0a0_20_0_fff;
invader_table[29]    <= 52'h8_090_0c0_20_0_fff;
invader_table[30]    <= 52'h8_090_0e0_20_0_fff;
invader_table[31]    <= 52'h8_090_100_20_0_fff;
invader_table[32]    <= 52'h0_020_1a0_20_0_fff;
invader_table[33]    <= 52'h0_020_1c0_20_0_fff;
invader_table[34]    <= 52'h0_020_1e0_20_0_fff;
invader_table[35]    <= 52'h0_020_200_20_0_fff;
invader_table[36]    <= 52'h0_020_220_20_0_fff;
invader_table[37]    <= 52'h0_020_240_20_0_fff;
invader_table[38]    <= 52'h0_020_260_20_0_fff;
invader_table[39]    <= 52'h0_000_000_20_0_000;
invader_table[40]    <= 52'h0_000_000_20_0_000;
invader_table[41]    <= 52'h0_000_000_20_0_000;
invader_table[42]    <= 52'h0_000_000_20_0_000;
invader_table[43]    <= 52'h0_000_000_20_0_000;
invader_table[44]    <= 52'h0_000_000_20_0_000;
invader_table[45]    <= 52'h0_000_000_20_0_000;
invader_table[46]    <= 52'h0_000_000_20_0_000;
invader_table[47]    <= 52'h0_000_000_20_0_000;
invader_table[48]    <= 52'h0_000_000_20_0_000;
invader_table[50]    <= 52'h0_1c0_000_20_1_fff;
invader_table[51]    <= 52'h0_000_000_20_0_000;
invader_table[52]    <= 52'h0_000_000_20_0_000;
invader_table[53]    <= 52'h0_000_000_20_0_000;
invader_table[54]    <= 52'h0_000_000_20_0_000;
invader_table[55]    <= 52'h0_000_000_20_0_000;
invader_table[56]    <= 52'h0_000_000_20_0_000;
invader_table[57]    <= 52'h0_000_000_20_0_000;
invader_table[58]    <= 52'h0_000_000_20_0_000;
invader_table[59]    <= 52'h0_000_000_20_0_000;
invader_table[60]    <= 52'h0_000_000_20_0_000;
invader_table[61]    <= 52'h0_1a0_000_20_1_000;
invader_table[62]    <= 52'h8_1c0_000_20_1_ff0;