                invT_pV[0] <= 8'h00;
                invT_pV[1] <= 8'h00;
                invT_pV[2] <= 8'h00;
                invT_pV[3] <= 8'h00;
                invT_pV[4] <= 8'h00;
                invT_pV[5] <= 8'h00;
                invT_pV[6] <= 8'h00;
                invT_pV[7] <= 8'h00;
                invT_pV[8] <= 8'h00;
                invT_pV[9] <= 8'h00;
                invT_pV[10] <= 8'h00;
                invT_pV[11] <= 8'h00;
                invT_pV[12] <= 8'h00;
                invT_pV[13] <= 8'h00;
                invT_pV[14] <= 8'h00;
                invT_pV[15] <= 8'h00;
                invT_pV[16] <= 8'h00;
                invT_pV[17] <= 8'h00;
                invT_pV[18] <= 8'h00;
                invT_pV[19] <= 8'h00;
                invT_pV[20] <= 8'h00;
                invT_pV[21] <= 8'h00;
                invT_pV[22] <= 8'h00;
                invT_pV[23] <= 8'h00;
                invT_pV[24] <= 8'h00;
                invT_pV[25] <= 8'h00;
                invT_pV[26] <= 8'h00;
                invT_pV[27] <= 8'h00;
                invT_pV[28] <= 8'h00;
                invT_pV[29] <= 8'h00;
                invT_pV[30] <= 8'h00;
                invT_pV[31] <= 8'h00;
                invT_pV[32] <= 8'h00;
                invT_pV[33] <= 8'h00;
                invT_pV[34] <= 8'h00;
                invT_pV[35] <= 8'h00;
                invT_pV[36] <= 8'h00;
                invT_pV[37] <= 8'h00;
                invT_pV[38] <= 8'h00;
                invT_pV[39] <= 8'h00;
                invT_pV[40] <= 8'h00;
                invT_pV[41] <= 8'h00;
                invT_pV[42] <= 8'h00;
                invT_pV[43] <= 8'h00;
                invT_pV[44] <= 8'h00;
                invT_pV[45] <= 8'h00;
                invT_pV[46] <= 8'h00;
                invT_pV[47] <= 8'h00;
                invT_pV[48] <= 8'h00;
                invT_pV[49] <= 8'h00;
                invT_pV[50] <= 8'h00;
                invT_pV[51] <= 8'h00;
                invT_pV[52] <= 8'h00;
                invT_pV[53] <= 8'h00;
                invT_pV[54] <= 8'h00;
                invT_pV[55] <= 8'h00;
                invT_pV[56] <= 8'h00;
                invT_pV[57] <= 8'h00;
                invT_pV[58] <= 8'h00;
                invT_pV[59] <= 8'h00;
                invT_pV[60] <= 8'h00;
                invT_pV[61] <= 8'h00;
                invT_pV[62] <= 8'h00;

                invT_pH[0] <= 8'h00;
                invT_pH[1] <= 8'h00;
                invT_pH[2] <= 8'h00;
                invT_pH[3] <= 8'h00;
                invT_pH[4] <= 8'h00;
                invT_pH[5] <= 8'h00;
                invT_pH[6] <= 8'h00;
                invT_pH[7] <= 8'h00;
                invT_pH[8] <= 8'h00;
                invT_pH[9] <= 8'h00;
                invT_pH[10] <= 8'h00;
                invT_pH[11] <= 8'h00;
                invT_pH[12] <= 8'h00;
                invT_pH[13] <= 8'h00;
                invT_pH[14] <= 8'h00;
                invT_pH[15] <= 8'h00;
                invT_pH[16] <= 8'h00;
                invT_pH[17] <= 8'h00;
                invT_pH[18] <= 8'h00;
                invT_pH[19] <= 8'h00;
                invT_pH[20] <= 8'h00;
                invT_pH[21] <= 8'h00;
                invT_pH[22] <= 8'h00;
                invT_pH[23] <= 8'h00;
                invT_pH[24] <= 8'h00;
                invT_pH[25] <= 8'h00;
                invT_pH[26] <= 8'h00;
                invT_pH[27] <= 8'h00;
                invT_pH[28] <= 8'h00;
                invT_pH[29] <= 8'h00;
                invT_pH[30] <= 8'h00;
                invT_pH[31] <= 8'h00;
                invT_pH[32] <= 8'h00;
                invT_pH[33] <= 8'h00;
                invT_pH[34] <= 8'h00;
                invT_pH[35] <= 8'h00;
                invT_pH[36] <= 8'h00;
                invT_pH[37] <= 8'h00;
                invT_pH[38] <= 8'h00;
                invT_pH[39] <= 8'h00;
                invT_pH[40] <= 8'h00;
                invT_pH[41] <= 8'h00;
                invT_pH[42] <= 8'h00;
                invT_pH[43] <= 8'h00;
                invT_pH[44] <= 8'h00;
                invT_pH[45] <= 8'h00;
                invT_pH[46] <= 8'h00;
                invT_pH[47] <= 8'h00;
                invT_pH[48] <= 8'h00;
                invT_pH[49] <= 8'h00;
                invT_pH[50] <= 8'h00;
                invT_pH[51] <= 8'h00;
                invT_pH[52] <= 8'h00;
                invT_pH[53] <= 8'h00;
                invT_pH[54] <= 8'h00;
                invT_pH[55] <= 8'h00;
                invT_pH[56] <= 8'h00;
                invT_pH[57] <= 8'h00;
                invT_pH[58] <= 8'h00;
                invT_pH[59] <= 8'h00;
                invT_pH[60] <= 8'h00;
                invT_pH[61] <= 8'h00;
                invT_pH[62] <= 8'h00;